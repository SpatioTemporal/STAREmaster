netcdf MOD05_L2.A2005349.2125.061.2017294065400_stare {
dimensions:
	i_5km = 406 ;
	j_5km = 270 ;
	l_5km = 7221 ;
variables:
	double Latitude_5km(i_5km, j_5km) ;
		Latitude_5km:long_name = "latitude" ;
		Latitude_5km:units = "degrees_north" ;
	double Longitude_5km(i_5km, j_5km) ;
		Longitude_5km:long_name = "longitude" ;
		Longitude_5km:units = "degrees_east" ;
	uint64 STARE_index_5km(i_5km, j_5km) ;
		STARE_index_5km:long_name = "SpatioTemporal Adaptive Resolution Encoding (STARE) index" ;
		STARE_index_5km:variables = "" ;
	uint64 STARE_cover_5km(l_5km) ;
		STARE_cover_5km:long_name = "SpatioTemporal Adaptive Resolution Encoding (STARE) cover" ;

// global attributes:
		:title = "SpatioTemporal Adaptive Resolution Encoding (STARE) sidecar file" ;
		:institution = "Institute for the Study of Institutes" ;
		:source = "STAREmaster 1.0.0" ;
}
